module Xor_gate(
	input a,b,
	output c
	);

xor xx1 (c,a,b);

endmodule
